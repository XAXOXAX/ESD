----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 16.11.2018 16:24:23
-- Design Name: 
-- Module Name: MUX - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MUX6b_01_12 is
  Port (    In1,In2: in std_logic_vector (5 downto 0);
            sel:in std_logic;
            SigOut: out std_logic_vector (5 downto 0));
end MUX6b_01_12;

architecture Behavioral of MUX6b_01_12 is

begin

SigOut<=In2 when (sel='1');
SigOut<=In1 when (sel='0');


end Behavioral;
